*** SPICE deck for cell tau_result{sch} from library to_calculate_cinv
*** Created on Mon May 03, 2021 23:11:11
*** Last revised on Sun May 16, 2021 13:58:50
*** Written on Sun May 16, 2021 13:59:43 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT to_calculate_cinv__inverter_size_1 FROM CELL inverter_size_1{sch}
.SUBCKT to_calculate_cinv__inverter_size_1 A F gnd vdd
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 F A gnd gnd N L=0.2U W=0.4U
Mpmos@0 vdd A F vdd P L=0.2U W=1U
.ENDS to_calculate_cinv__inverter_size_1

.global gnd vdd

*** TOP LEVEL CELL: tau_result{sch}
Rres@0 out in 10k
Xinverter@0 out f gnd vdd to_calculate_cinv__inverter_size_1

* Spice Code nodes in cell cell 'tau_result{sch}'
vdd vdd 0 dc 1.8
vin in 0 pulse 0 1.8 10n 0p 0p 20n 50n
.measure tau trig v(out) val=0 rise=1 TARG v(out) val=1.1376 rise=1
.tran 0 200n
.include D:\AUC\8th Semester - Spring 21\DD2\Project\scmos18.txt
.END
